module Reg(Clk, RegWr, busW, Rw, Ra, Rb, busA, busB);
// ���룺ʱ���ź�,�Ĵ���дʹ���ź�,�Ĵ���д������,��ȡ����A,��ȡ����B,д������
// ��������A,���B

	input Clk, RegWr, Rw, Ra, Rb, busW;

	output reg [31:0] busA, busB;

	//parameter n = 32; // �Ĵ���λ��

	reg [31:0] regs[31:0]; // 32��32λ�Ĵ���������

	integer i;

	initial begin
		// ��ʼ���Ĵ��������ǰ����Ԫ��
		regs[0] = 32'h00000000;
		regs[1] = 32'h00000012; // 18
		regs[2] = 32'h00000024; // 36
		regs[3] = 32'h00000102; // 258
		regs[4] = 32'h00000063; // 99
		// ������Ԫ�س�ʼ��Ϊ0
		for (i = 5; i < 32; i = i + 1) regs[i] = 32'h0;
	end

	// дʹ���ź���Чʱ��д������д��ָ���Ĵ���
	always @(negedge Clk) begin
		if (RegWr == 1) regs[Rw] <= busW;
	end

	// ����ȡ�Ĵ���A��B�����������仯ʱ���ӼĴ��������ж�ȡ��Ӧ�����ݲ������������
	always @(Ra or Rb) begin
		busA <= regs[Ra];
		busB <= regs[Rb];
	end
endmodule
